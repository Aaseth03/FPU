LIBRARY ieee;
USE ieee.STD_LOGIC_1164.all;
USE ieee.STD_LOGIC_UNSIGNED.all;
USE ieee.NUMERIC_STD.all;
-- Teller antall 0'er før ledende 1'er
ENTITY Z_COUNTER IS
	PORT(
		addresult	:	IN		UNSIGNED(24 DOWNTO 0);
		Zeros			:	OUT	NATURAL := 0
		);
END Z_COUNTER;

ARCHITECTURE Struct OF Z_COUNTER IS
	SIGNAL	b24,b23,b22,b21,b20,b19,b18,b17,b16,b15,b14,b13,b12,b11,b10,b9,b8,b7,b6,b5,b4,b3,b2,b1,b0 : NATURAL RANGE 0 to 1 := 0;
	SIGNAL	tmp	:	UNSIGNED(24 DOWNTO 0);
BEGIN
	
	tmp <= NOT(addresult);
	
	PROCESS(tmp, b24,b23,b22,b21,b20,b19,b18,b17,b16,b15,b14,b13,b12,b11,b10,b9,b8,b7,b6,b5,b4,b3,b2,b1,b0)
	BEGIN
		IF((tmp AND ("1000000000000000000000000")) = "1000000000000000000000000") THEN
			b24 <= 1;
		ELSE
			b24 <= 0;
		END IF;
		IF((tmp AND ("1100000000000000000000000")) = "1100000000000000000000000") THEN
			b23 <= 1;
		ELSE
			b23 <= 0;
		END IF;
		IF((tmp AND ("1110000000000000000000000")) = "1110000000000000000000000") THEN
			b22 <= 1;
		ELSE
			b22 <= 0;
		END IF;
		IF((tmp AND ("1111000000000000000000000")) = "1111000000000000000000000") THEN
			b21 <= 1;
		ELSE
			b21 <= 0;
		END IF;
		IF((tmp AND ("1111100000000000000000000")) = "1111100000000000000000000") THEN
			b20 <= 1;
		ELSE
			b20 <= 0;
		END IF;
		IF((tmp AND ("1111110000000000000000000")) = "1111110000000000000000000") THEN
			b19 <= 1;
		ELSE
			b19 <= 0;
		END IF;
		IF((tmp AND ("1111111000000000000000000")) = "1111111000000000000000000") THEN
			b18 <= 1;
		ELSE
			b18 <= 0;
		END IF;
		IF((tmp AND ("1111111100000000000000000")) = "1111111100000000000000000") THEN
			b17 <= 1;
		ELSE
			b17 <= 0;
		END IF;
		IF((tmp AND ("1111111110000000000000000")) = "1111111110000000000000000") THEN
			b16 <= 1;
		ELSE
			b16 <= 0;
		END IF;
		IF((tmp AND ("1111111111000000000000000")) = "1111111111000000000000000") THEN
			b15 <= 1;
		ELSE
			b15 <= 0;
		END IF;
		IF((tmp AND ("1111111111100000000000000")) = "1111111111100000000000000") THEN
			b14 <= 1;
		ELSE
			b14 <= 0;
		END IF;
		IF((tmp AND ("1111111111110000000000000")) = "1111111111110000000000000") THEN
			b13 <= 1;
		ELSE
			b13 <= 0;
		END IF;
		IF((tmp AND ("1111111111111000000000000")) = "1111111111111000000000000") THEN
			b12 <= 1;
		ELSE
			b12 <= 0;
		END IF;
		IF((tmp AND ("1111111111111100000000000")) = "1111111111111100000000000") THEN
			b11 <= 1;
		ELSE
			b11 <= 0;
		END IF;
		IF((tmp AND ("1111111111111110000000000")) = "1111111111111110000000000") THEN
			b10 <= 1;
		ELSE
			b10 <= 0;
		END IF;
		IF((tmp AND ("1111111111111111000000000")) = "1111111111111111000000000") THEN
			b9 <= 1;
		ELSE
			b9 <= 0;
		END IF;
		IF((tmp AND ("1111111111111111100000000")) = "1111111111111111100000000") THEN
			b8 <= 1;
		ELSE
			b8 <= 0;
		END IF;
		IF((tmp AND ("1111111111111111110000000")) = "1111111111111111110000000") THEN
			b7 <= 1;
		ELSE
			b7 <= 0;
		END IF;
		IF((tmp AND ("1111111111111111111000000")) = "1111111111111111111000000") THEN
			b6 <= 1;
		ELSE
			b6 <= 0;
		END IF;
		IF((tmp AND ("1111111111111111111100000")) = "1111111111111111111100000") THEN
			b5 <= 1;
		ELSE
			b5 <= 0;
		END IF;
		IF((tmp AND ("1111111111111111111110000")) = "1111111111111111111110000") THEN
			b4 <= 1;
		ELSE
			b4 <= 0;
		END IF;
		IF((tmp AND ("1111111111111111111111000")) = "1111111111111111111111000") THEN
			b3 <= 1;
		ELSE
			b3 <= 0;
		END IF;
		IF((tmp AND ("1111111111111111111111100")) = "1111111111111111111111100") THEN
			b2 <= 1;
		ELSE
			b2 <= 0;
		END IF;
		IF((tmp AND ("1111111111111111111111110")) = "1111111111111111111111110") THEN
			b1 <= 1;
		ELSE
			b1 <= 0;
		END IF;
		IF((tmp AND ("1111111111111111111111111")) = "1111111111111111111111111") THEN
			b0 <= 1;
		ELSE
			b0 <= 0;
		END IF;
		Zeros <= (b24+b23+b22+b21+b20+b19+b18+b17+b16+b15+b14+b13+b12+b11+b10+b9+b8+b7+b6+b5+b4+b3+b2+b1+b0);

	END PROCESS;
END Struct;



	